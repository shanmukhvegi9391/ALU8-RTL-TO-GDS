VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu8
  CLASS BLOCK ;
  FOREIGN alu8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.670 BY 81.390 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 68.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 68.240 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 66.670 17.040 70.670 17.640 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 66.670 20.440 70.670 21.040 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 77.390 26.130 81.390 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 77.390 42.230 81.390 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 66.670 47.640 70.670 48.240 ;
    END
  END b[7]
  PIN carry_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 66.670 54.440 70.670 55.040 ;
    END
  END carry_out
  PIN negative
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 77.390 51.890 81.390 ;
    END
  END negative
  PIN op[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 66.670 44.240 70.670 44.840 ;
    END
  END op[0]
  PIN op[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 66.670 37.440 70.670 38.040 ;
    END
  END op[1]
  PIN op[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 66.670 40.840 70.670 41.440 ;
    END
  END op[2]
  PIN op[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 66.670 34.040 70.670 34.640 ;
    END
  END op[3]
  PIN overflow
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 66.670 57.840 70.670 58.440 ;
    END
  END overflow
  PIN y[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 77.390 39.010 81.390 ;
    END
  END y[0]
  PIN y[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END y[2]
  PIN y[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END y[3]
  PIN y[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END y[4]
  PIN y[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 77.390 32.570 81.390 ;
    END
  END y[5]
  PIN y[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 77.390 35.790 81.390 ;
    END
  END y[6]
  PIN y[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 77.390 48.670 81.390 ;
    END
  END y[7]
  PIN zero
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 77.390 45.450 81.390 ;
    END
  END zero
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 65.050 68.190 ;
      LAYER li1 ;
        RECT 5.520 10.795 64.860 68.085 ;
      LAYER met1 ;
        RECT 4.210 10.640 64.860 68.240 ;
      LAYER met2 ;
        RECT 4.230 77.110 25.570 77.930 ;
        RECT 26.410 77.110 32.010 77.930 ;
        RECT 32.850 77.110 35.230 77.930 ;
        RECT 36.070 77.110 38.450 77.930 ;
        RECT 39.290 77.110 41.670 77.930 ;
        RECT 42.510 77.110 44.890 77.930 ;
        RECT 45.730 77.110 48.110 77.930 ;
        RECT 48.950 77.110 51.330 77.930 ;
        RECT 52.170 77.110 63.850 77.930 ;
        RECT 4.230 4.280 63.850 77.110 ;
        RECT 4.230 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 63.850 4.280 ;
      LAYER met3 ;
        RECT 3.990 58.840 66.670 68.165 ;
        RECT 3.990 57.440 66.270 58.840 ;
        RECT 3.990 55.440 66.670 57.440 ;
        RECT 4.400 54.040 66.270 55.440 ;
        RECT 3.990 52.040 66.670 54.040 ;
        RECT 4.400 50.640 66.670 52.040 ;
        RECT 3.990 48.640 66.670 50.640 ;
        RECT 4.400 47.240 66.270 48.640 ;
        RECT 3.990 45.240 66.670 47.240 ;
        RECT 4.400 43.840 66.270 45.240 ;
        RECT 3.990 41.840 66.670 43.840 ;
        RECT 4.400 40.440 66.270 41.840 ;
        RECT 3.990 38.440 66.670 40.440 ;
        RECT 4.400 37.040 66.270 38.440 ;
        RECT 3.990 35.040 66.670 37.040 ;
        RECT 4.400 33.640 66.270 35.040 ;
        RECT 3.990 31.640 66.670 33.640 ;
        RECT 4.400 30.240 66.670 31.640 ;
        RECT 3.990 28.240 66.670 30.240 ;
        RECT 4.400 26.840 66.670 28.240 ;
        RECT 3.990 21.440 66.670 26.840 ;
        RECT 3.990 20.040 66.270 21.440 ;
        RECT 3.990 18.040 66.670 20.040 ;
        RECT 3.990 16.640 66.270 18.040 ;
        RECT 3.990 10.715 66.670 16.640 ;
      LAYER met4 ;
        RECT 17.775 17.855 20.640 58.305 ;
        RECT 23.040 17.855 23.940 58.305 ;
        RECT 26.340 17.855 47.545 58.305 ;
  END
END alu8
END LIBRARY

